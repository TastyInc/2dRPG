? %)': $s<-25$!<. lps}ak|qstqcl1?-86>2'-5 lpc|ab|qs}qclps<-25$!%56!2s}aalrsxaflw
savefile playerpos 1 1 800 800 playerstats 100 100 100 1 playeritems 1 2 3 4 5 6