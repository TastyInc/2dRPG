savefile playerpos 1 1 453 150 playerstats 100 100 100 1 playeritems 1 2 3 4 5 666