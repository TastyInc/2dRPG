playerpos maptheme mapscreen x y
playerstats health endurance strenght dexterity oder so
playeritems gun sword angere shit
gametime time